-- SPDX-License-Identifier: MIT
-- Copyright (c) 2021 Ross K. Snider.  All rights reserved.
----------------------------------------------------------------------------
-- Description:  Template for Synchronous VHDL Process
----------------------------------------------------------------------------
-- Author:       Ross K. Snider
-- Company:      Montana State University
-- Create Date:  September 30, 2021
-- Revision:     1.0
-- License: MIT  (opensource.org/licenses/MIT)
----------------------------------------------------------------------------

my_synchronous_process : process(clk)
begin
    if rising_edge(clk) then 
	 
        -- insert synchronous logic here
		  
    end if;
end process;
