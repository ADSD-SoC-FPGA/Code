
add code 
